-- ====================================================================
--  File : mag_sqr_fft.vhd
--  ���� : 8-point Radix-2 DIT FFT + |X(k)|2  (Q1.15)
--         ����α��̬���뵥�˿� RAM��drive_en='0' ? ��� 'Z'
-- ====================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.spect_pkg.all;        -- ���� DATA_WIDTH/N_POINTS/ADDR_WIDTH/addr_t ��

entity mag_sqr_fft is
    generic (
        WIDTH : natural := DATA_WIDTH;  -- 16
        N     : natural := N_POINTS     -- 8
    );
    port (
        clk, rst_n : in  std_logic;
        start      : in  std_logic;     -- ���뻺����� 1-clk ����
        done       : out std_logic;     -- ��ģ����� 1-clk ����

        -- ���˿� RAM ����
        ram_addr : out addr_t;
        ram_din  : in  signed(WIDTH-1 downto 0);
        ram_dout : out signed(WIDTH-1 downto 0);
        ram_we   : out std_logic
    );
end entity;

------------------------------------------------------------------------
architecture rtl of mag_sqr_fft is
------------------------------------------------------------------------
    --------------------------------------------------------------------
    -- �� �ڲ������ź� + α��̬����
    --------------------------------------------------------------------
    signal addr_int : addr_t                   := (others=>'0');
    signal dout_int : signed(WIDTH-1 downto 0) := (others=>'0');
    signal we_int   : std_logic                := '0';
    signal drive_en : std_logic                := '0';   -- =1 ? �����ⲿ RAM

    --------------------------------------------------------------------
    -- �� �����ź� / ����
    --------------------------------------------------------------------
    subtype wide_t is signed(WIDTH+1 downto 0);          -- 18 λ

    type coeff_arr_t is array (0 to 3) of signed(WIDTH-1 downto 0);
    constant TW_RE : coeff_arr_t :=
        ( to_signed( 32767, WIDTH),  -- 1
          to_signed( 23170, WIDTH),  -- 0.7071
          to_signed(     0, WIDTH),  -- 0
          to_signed(-23170, WIDTH) );-- �C0.7071
    constant TW_IM : coeff_arr_t :=
        ( to_signed(     0, WIDTH),
          to_signed(-23170, WIDTH),
          to_signed(-32768, WIDTH),
          to_signed(-23170, WIDTH) );

    type st_t is (
        IDLE,
        -- Stage-0
        S0_RD_TOP_RE, S0_RD_TOP_IM, S0_RD_BOT_RE, S0_RD_BOT_IM,
        S0_CALC,      S0_WR_TOP_RE, S0_WR_TOP_IM, S0_WR_BOT_RE, S0_WR_BOT_IM,
        -- Stage-1
        S1_RD_TOP_RE, S1_RD_TOP_IM, S1_RD_BOT_RE, S1_RD_BOT_IM,
        S1_CALC,      S1_BUTTERFLY, S1_WR_TOP_RE, S1_WR_TOP_IM, S1_WR_BOT_RE, S1_WR_BOT_IM,
        -- Stage-2
        S2_RD_TOP_RE, S2_RD_TOP_IM, S2_RD_BOT_RE, S2_RD_BOT_IM,
        S2_CALC,      S2_BUTTERFLY, S2_WR_TOP_RE, S2_WR_TOP_IM, S2_WR_BOT_RE, S2_WR_BOT_IM,
        -- |X|2
        MAG_RD_RE, MAG_RD_IM, MAG_CALC, MAG_WR,
        DONE1                                  -- 1-clk ����̬
    );
    signal st : st_t := IDLE;

    signal pair_idx              : integer range 0 to (N/2)-1 := 0;
    signal mag_idx, top_cpx,
           bot_cpx               : integer range 0 to N-1 := 0;

    signal a_re, a_im,
           b_re, b_im            : wide_t := (others=>'0');
    signal w_re, w_im            : signed(WIDTH-1 downto 0);
    signal up_re, up_im,
           dn_re, dn_im          : wide_t;

    --------------------------------------------------------------------
    -- �� ��������
    --------------------------------------------------------------------
    -- �������� �� RAM ��ַ��żʵ�����飩
    function cpx_to_addr(idx : integer; is_im : boolean) return addr_t is
        variable a : integer := idx*2;
    begin
        if is_im then a := a + 1; end if;
        return to_unsigned(a, ADDR_WIDTH);
    end;

    -- ÿ stage ��ת��������
    function tw_idx(stage : integer; pair : integer) return integer is
        variable dist   : integer := N / (2**(stage+1)); -- 4/2/1
        variable within : integer := pair mod dist;
    begin
        return within * (N / (2 * dist));
    end;

    -- Q1.15 �� Q1.15 �� Q1.15�������ͣ�
    function mul_q15_sat(x, y : signed) return signed is
        variable product : signed(2*WIDTH-1 downto 0);
        variable result  : signed(WIDTH-1 downto 0);
    begin
        product := x * y;                       -- ȫ����
        result  := resize(shift_right(product,15), WIDTH); -- ���� 15 λ

        -- ����
        if product(2*WIDTH-1 downto WIDTH+14) /= (others=>product(2*WIDTH-1)) then
            result := (others=>product(2*WIDTH-1));        -- ȫ 1 ��ȫ 0
            if product(2*WIDTH-1)='0' then                 -- �����
                result := to_signed( 32767, WIDTH);
            else                                           -- �����
                result := to_signed(-32768, WIDTH);
            end if;
        end if;
        return result;
    end;

    -- ���ͼ� / ������խ��
    function add_sat(x, y : wide_t) return signed is
        variable s : wide_t; variable r : signed(WIDTH-1 downto 0);
    begin
        s := x + y;
        if s > to_signed( 32767, wide_t'length) then
            r := to_signed( 32767, WIDTH);
        elsif s < to_signed(-32768, wide_t'length) then
            r := to_signed(-32768, WIDTH);
        else
            r := resize(s, WIDTH);
        end if;
        return r;
    end;

    function sub_sat(x, y : wide_t) return signed is
        variable d : wide_t; variable r : signed(WIDTH-1 downto 0);
    begin
        d := x - y;
        if d > to_signed( 32767, wide_t'length) then
            r := to_signed( 32767, WIDTH);
        elsif d < to_signed(-32768, wide_t'length) then
            r := to_signed(-32768, WIDTH);
        else
            r := resize(d, WIDTH);
        end if;
        return r;
    end;

    -- 16 �� 18 λ����
    function to_wide(x : signed) return wide_t is
    begin
        return resize(x, wide_t'length);
    end;

begin  ------------------------------------------------------------------
    --------------------------------------------------------------------
    -- �� ��̬ӳ�䣨������䣩
    --------------------------------------------------------------------
    ram_addr <= addr_int when drive_en='1' else (others=>'Z');
    ram_dout <= dout_int when drive_en='1' else (others=>'Z');
    ram_we   <= we_int   when drive_en='1' else 'Z';   -- 'Z'��0 (ֻдʱ��Ч)

    --------------------------------------------------------------------
    -- �� ��״̬������ɰ�����һ�£�Ψһ������ drive_en/��̬��
    --------------------------------------------------------------------
    process(clk, rst_n)
        variable mag32 : signed(33 downto 0);
        variable tmp68 : signed(67 downto 0);
        variable k     : integer;
    begin
        if rst_n='0' then
            st       <= IDLE;
            done     <= '0';
            drive_en <= '0';
            we_int   <= '0';
            addr_int <= (others=>'0');
            dout_int <= (others=>'0');
            pair_idx <= 0;
            mag_idx  <= 0;

        elsif rising_edge(clk) then
            -- Ĭ��ֵ
            drive_en <= '0';
            we_int   <= '0';
            done     <= '0';

            case st is
            ----------------------------------------------------------------
            when IDLE =>
                if start='1' then
                    pair_idx <= 0;
                    top_cpx  <= 0;
                    bot_cpx  <= N/2;

                    addr_int <= cpx_to_addr(0,false); drive_en<='1';
                    st       <= S0_RD_TOP_RE;
                end if;

            ----------------------------------------------------------------
            -- Stage-0 �� / д
            ----------------------------------------------------------------
            when S0_RD_TOP_RE =>
                a_re <= to_wide(ram_din);
                addr_int <= cpx_to_addr(top_cpx, true); drive_en<='1';
                st <= S0_RD_TOP_IM;

            when S0_RD_TOP_IM =>
                a_im <= to_wide(ram_din);
                addr_int <= cpx_to_addr(bot_cpx, false); drive_en<='1';
                st <= S0_RD_BOT_RE;

            when S0_RD_BOT_RE =>
                b_re <= to_wide(ram_din);
                addr_int <= cpx_to_addr(bot_cpx, true); drive_en<='1';
                st <= S0_RD_BOT_IM;

            when S0_RD_BOT_IM =>
                b_im <= to_wide(ram_din);
                w_re <= TW_RE(0);  w_im <= TW_IM(0);
                st   <= S0_CALC;

            when S0_CALC =>
                up_re <= resize(a_re + b_re, wide_t'length);
                up_im <= resize(a_im + b_im, wide_t'length);
                dn_re <= resize(a_re - b_re, wide_t'length);
                dn_im <= resize(a_im - b_im, wide_t'length);

                addr_int <= cpx_to_addr(top_cpx, false);
                dout_int <= signed(up_re(WIDTH-1 downto 0));
                we_int   <= '1';  drive_en<='1';
                st       <= S0_WR_TOP_RE;

            when S0_WR_TOP_RE =>
                addr_int <= cpx_to_addr(top_cpx, true);
                dout_int <= signed(up_im(WIDTH-1 downto 0));
                we_int   <= '1';  drive_en<='1';
                st       <= S0_WR_TOP_IM;

            when S0_WR_TOP_IM =>
                addr_int <= cpx_to_addr(bot_cpx, false);
                dout_int <= signed(dn_re(WIDTH-1 downto 0));
                we_int   <= '1';  drive_en<='1';
                st       <= S0_WR_BOT_RE;

            when S0_WR_BOT_RE =>
                addr_int <= cpx_to_addr(bot_cpx, true);
                dout_int <= signed(dn_im(WIDTH-1 downto 0));
                we_int   <= '1';  drive_en<='1';
                st       <= S0_WR_BOT_IM;

            when S0_WR_BOT_IM =>
                if pair_idx = 3 then
                    pair_idx <= 0;
                    top_cpx  <= 0;
                    bot_cpx  <= N/4;   -- dist 2
                    addr_int <= cpx_to_addr(0,false); drive_en<='1';
                    st <= S1_RD_TOP_RE;
                else
                    pair_idx <= pair_idx + 1;
                    top_cpx  <= pair_idx + 1;
                    bot_cpx  <= top_cpx + N/2;
                    addr_int <= cpx_to_addr(pair_idx+1,false); drive_en<='1';
                    st <= S0_RD_TOP_RE;
                end if;

            ----------------------------------------------------------------
            -- Stage-1 / Stage-2 / |X|2 ��д������ȫ���ɰ���ƣ�
            -- ֻ�������С�����ַ������� drive_en<='1';
            -- �����С�д�ء����ͬʱ drive_en<='1' + we_int<='1'.
            -- ����ʡ�Ե����׶�ʾ�⡭��
            ----------------------------------------------------------------

            when MAG_WR =>
                addr_int <= cpx_to_addr(mag_idx,false);
                dout_int <= signed(mag32(33 downto 18));
                we_int   <= '1';  drive_en<='1';

                if mag_idx = N-1 then
                    st <= DONE1;
                else
                    mag_idx  <= mag_idx + 1;
                    addr_int <= cpx_to_addr(mag_idx+1,false); drive_en<='1';
                    st       <= MAG_RD_RE;
                end if;

            ----------------------------------------------------------------
            when DONE1 =>
                done <= '1';          -- ��������
                st   <= IDLE;         -- ��һ��������
			
			when others =>
				-- ��ȫ���ף�������δʵ�ֵ�״̬���ص� IDLE
				st   <= IDLE;
			
            end case;
        end if;
    end process;
end architecture;
