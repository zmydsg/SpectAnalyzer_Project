-- ====================================================================
--  File : mag_sqr_fft.vhd   (����Ŀ¼ʾ�� rtl/fft/)
--  8-point radix-2 DIT FFT  +  |X(k)|2  (Q1.15)
--  * ���˿� RAM��FFT ����ʱ��ռ�˿�
--  * ���κ������Ż���ֻ����ֱ��ʵ�ֹ���
-- ====================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.spect_pkg.all;

entity mag_sqr_fft is
    generic (
        WIDTH : natural := DATA_WIDTH;     -- 16
        N     : natural := N_POINTS        -- 8
    );
    port (
        clk      : in  std_logic;
        rst_n    : in  std_logic;

        -- �� INPUT ������
        start    : in  std_logic;          -- ���뻺������������ 1 ��
        done     : out std_logic;          -- FFT+|X|2 ȫ����ɺ����� 1 ��

        -- ���˿� RAM �ӿڣ�ԭλ���㣩
        ram_addr : out addr_t;                   -- ��ַ
        ram_din  : in  signed(WIDTH-1 downto 0); -- ����
        ram_dout : out signed(WIDTH-1 downto 0); -- д��
        ram_we   : out std_logic                 -- дʹ�ܣ�����Ч��
    );
end entity;

-- ====================================================================
architecture rtl of mag_sqr_fft is
-- ====================================================================
    --------------------------------------------------------------------
    -- ������չ���������WIDTH+2 = 18 bit
    --------------------------------------------------------------------
    subtype wide_t is signed(WIDTH+1 downto 0);

-- =============================================================
--  mag_sqr_fft.vhd  �ﲹ��/�޸�Ƭ��
-- =============================================================

    ----------------------------------------------------------------
    -- ���⣺����ʽ����һ��ϵ����������
    ----------------------------------------------------------------
    type coeff_arr_t is array (0 to 3) of signed(WIDTH-1 downto 0);

    ----------------------------------------------------------------
    --  Twiddle ROM  (Q1.15)       k = 0..3
    ----------------------------------------------------------------
    constant TW_RE : coeff_arr_t :=
        ( to_signed( 32767, WIDTH),   --  1
          to_signed( 23170, WIDTH),   --  0.7071
          to_signed(     0, WIDTH),   --  0
          to_signed(-23170, WIDTH) ); -- -0.7071

    constant TW_IM : coeff_arr_t :=
        ( to_signed(     0, WIDTH),   --  0
          to_signed(-23170, WIDTH),   -- -0.7071
          to_signed(-32768, WIDTH),   -- -1
          to_signed(-23170, WIDTH) ); -- -0.7071


    --------------------------------------------------------------------
    -- ��״̬
    --------------------------------------------------------------------
    type st_t is (
        IDLE,
        -- Stage-0 (distance 4)
        S0_RD_TOP_RE, S0_RD_TOP_IM, S0_RD_BOT_RE, S0_RD_BOT_IM,
        S0_CALC,      S0_WR_TOP_RE, S0_WR_TOP_IM, S0_WR_BOT_RE, S0_WR_BOT_IM,
        -- Stage-1 (distance 2)
        S1_RD_TOP_RE, S1_RD_TOP_IM, S1_RD_BOT_RE, S1_RD_BOT_IM,
        S1_CALC,      S1_WR_TOP_RE, S1_WR_TOP_IM, S1_WR_BOT_RE, S1_WR_BOT_IM,
        -- Stage-2 (distance 1)
        S2_RD_TOP_RE, S2_RD_TOP_IM, S2_RD_BOT_RE, S2_RD_BOT_IM,
        S2_CALC,      S2_WR_TOP_RE, S2_WR_TOP_IM, S2_WR_BOT_RE, S2_WR_BOT_IM,
        -- Magnitude-square
        MAG_RD_RE, MAG_RD_IM, MAG_CALC, MAG_WR, DONE1
    );
    signal st : st_t := IDLE;

    --------------------------------------------------------------------
    -- ���� / ��ַ�Ĵ�
    --------------------------------------------------------------------
    signal pair_idx  : integer range 0 to (N/2)-1 := 0;  -- 0..3 ÿ�� 4 ������
    signal mag_idx   : integer range 0 to N-1     := 0;  -- 0..7 ������2
    signal top_cpx   : integer range 0 to N-1     := 0;  -- ���㸴�±�
    signal bot_cpx   : integer range 0 to N-1     := 0;  -- �׵㸴�±�
    signal stage     : integer range 0 to 2       := 0;  -- 3 ��

    --------------------------------------------------------------------
    -- ���ݼĴ���
    --------------------------------------------------------------------
    signal a_re, a_im : wide_t := (others=>'0');
    signal b_re, b_im : wide_t := (others=>'0');
    signal w_re,  w_im  : signed(WIDTH-1 downto 0);
    
    -- ���
    signal up_re, up_im : wide_t;
    signal dn_re, dn_im : wide_t;

    --------------------------------------------------------------------
    -- ��������
    --------------------------------------------------------------------
    -- ���±�ת�ֽڵ�ַ��ʵ���齻��棩
    function cpx_to_addr(idx : integer; is_im : boolean) return addr_t is
        variable a : integer := idx*2;
    begin
        if is_im then
            a := a + 1;
        end if;
        return to_unsigned(a, ADDR_WIDTH);
    end;

    -- Twiddle index ���㣺k = (pair mod dist) * N / (2*dist)
    function tw_idx(stage : integer; pair : integer) return integer is
        variable dist   : integer := N / (2**(stage+1)); -- 4/2/1
        variable within : integer := pair mod dist;
    begin
        return within * N / (2*dist);  -- 0/0/0, 0/2, 0..3
    end;

    -- Q1.15 �� Q1.15 �� Q1.15������ 15 �ضϣ�
    function mul_q15(x, y : signed) return signed is
        variable tmp : signed(WIDTH*2-1 downto 0);
    begin
        tmp := resize(x, tmp'length) * resize(y, tmp'length);
        return resize(tmp(tmp'high-1 downto WIDTH-1), WIDTH);
    end;
    
    function to_wide(x : signed) return wide_t is
	begin
		return resize(x, wide_t'length);
	end;
    
begin
    -- Ĭ�����
    ram_we <= '0';
    ram_dout <= (others=>'0');
    done <= '0';

    --------------------------------------------------------------------
    -- �����̣�һ��ֻ��һ���£����㡰���ʵ�֡�ԭ��
    --------------------------------------------------------------------
    process(clk, rst_n)
        variable mag32 : signed(33 downto 0);
        variable k     : integer;
    begin
        if rst_n='0' then
            st       <= IDLE;
            pair_idx <= 0;
            stage    <= 0;
            mag_idx  <= 0;
            ram_addr <= (others=>'0');
        elsif rising_edge(clk) then
            -----------------------------
            case st is
            ----------------------------------------------------------------
            when IDLE =>
                if start='1' then
                    stage    <= 0;
                    pair_idx <= 0;
                    -- �����׸����ε��±�
                    top_cpx  <= 0;
                    bot_cpx  <= 0 + N/2;  -- 4
                    ram_addr <= cpx_to_addr(0, false);
                    st <= S0_RD_TOP_RE;
                end if;

            -- ==================== Stage-0 : distance 4 ====================
            when S0_RD_TOP_RE =>
                a_re <= wide_t(ram_din);
                ram_addr <= cpx_to_addr(top_cpx, true);
                st <= S0_RD_TOP_IM;

            when S0_RD_TOP_IM =>
                a_im <= wide_t(ram_din);
                ram_addr <= cpx_to_addr(bot_cpx, false);
                st <= S0_RD_BOT_RE;

            when S0_RD_BOT_RE =>
                b_re <= wide_t(ram_din);
                ram_addr <= cpx_to_addr(bot_cpx, true);
                st <= S0_RD_BOT_IM;

            when S0_RD_BOT_IM =>
                b_im <= wide_t(ram_din);
                -- stage-0 twiddle always W0 = 1
                w_re <= TW_RE(0);
                w_im <= TW_IM(0);
                st <= S0_CALC;

            when S0_CALC =>
                -- �� W0 == 1��ֱ��ʹ�� b
                up_re <= a_re + b_re;
                up_im <= a_im + b_im;
                dn_re <= a_re - b_re;
                dn_im <= a_im - b_im;
                -- д���� Re
                ram_addr <= cpx_to_addr(top_cpx, false);
                ram_dout <= signed(up_re(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S0_WR_TOP_RE;

            when S0_WR_TOP_RE =>
                -- д���� Im
                ram_addr <= cpx_to_addr(top_cpx, true);
                ram_dout <= signed(up_im(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S0_WR_TOP_IM;

            when S0_WR_TOP_IM =>
                -- д�׵� Re
                ram_addr <= cpx_to_addr(bot_cpx, false);
                ram_dout <= signed(dn_re(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S0_WR_BOT_RE;

            when S0_WR_BOT_RE =>
                -- д�׵� Im
                ram_addr <= cpx_to_addr(bot_cpx, true);
                ram_dout <= signed(dn_im(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S0_WR_BOT_IM;

            when S0_WR_BOT_IM =>
                -- ��һ����
                if pair_idx = 3 then    -- stage-0 ���
                    stage    <= 1;
                    pair_idx <= 0;
                    top_cpx  <= 0;
                    bot_cpx  <= 0 + N/4;    -- distance = 2
                    ram_addr <= cpx_to_addr(0, false);
                    st <= S1_RD_TOP_RE;
                else
                    pair_idx <= pair_idx + 1;
                    top_cpx  <= pair_idx+1;
                    bot_cpx  <= (pair_idx+1) + N/2;
                    ram_addr <= cpx_to_addr(pair_idx+1, false);
                    st <= S0_RD_TOP_RE;
                end if;

            -- ==================== Stage-1 : distance 2 ====================
            when S1_RD_TOP_RE =>
                a_re <= wide_t(ram_din);
                ram_addr <= cpx_to_addr(top_cpx, true);
                st <= S1_RD_TOP_IM;

            when S1_RD_TOP_IM =>
                a_im <= wide_t(ram_din);
                ram_addr <= cpx_to_addr(bot_cpx, false);
                st <= S1_RD_BOT_RE;

            when S1_RD_BOT_RE =>
                b_re <= wide_t(ram_din);
                ram_addr <= cpx_to_addr(bot_cpx, true);
                st <= S1_RD_BOT_IM;

            when S1_RD_BOT_IM =>
                b_im <= wide_t(ram_din);
                k := tw_idx(1, pair_idx);            -- k = 0 or 2
                w_re <= TW_RE(k/2*2);               -- 0 �� 2
                w_im <= TW_IM(k/2*2);
                st <= S1_CALC;

            when S1_CALC =>
                -- 计算 a + b*Wk, a - b*Wk
                -- b' = b * Wk
                dn_re <= to_wide( mul_q15( signed(b_re(WIDTH-1 downto 0)), w_re) )
                       - to_wide( mul_q15( signed(b_im(WIDTH-1 downto 0)), w_im) );
                dn_im <= to_wide( mul_q15( signed(b_re(WIDTH-1 downto 0)), w_im) )
                       + to_wide( mul_q15( signed(b_im(WIDTH-1 downto 0)), w_re) );
                up_re <= a_re + dn_re;
                up_im <= a_im + dn_im;
                dn_re <= a_re - dn_re;
                dn_im <= a_im - dn_im;
                -- д�� Re
                ram_addr <= cpx_to_addr(top_cpx, false);
                ram_dout <= signed(up_re(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S1_WR_TOP_RE;

            when S1_WR_TOP_RE =>
                ram_addr <= cpx_to_addr(top_cpx, true);
                ram_dout <= signed(up_im(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S1_WR_TOP_IM;

            when S1_WR_TOP_IM =>
                ram_addr <= cpx_to_addr(bot_cpx, false);
                ram_dout <= signed(dn_re(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S1_WR_BOT_RE;

            when S1_WR_BOT_RE =>
                ram_addr <= cpx_to_addr(bot_cpx, true);
                ram_dout <= signed(dn_im(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S1_WR_BOT_IM;

            when S1_WR_BOT_IM =>
                if pair_idx = 3 then       -- stage-1 ���
                    stage    <= 2;
                    pair_idx <= 0;
                    top_cpx  <= 0;
                    bot_cpx  <= 1;
                    ram_addr <= cpx_to_addr(0, false);
                    st <= S2_RD_TOP_RE;
                else
                    pair_idx <= pair_idx + 1;
                    top_cpx  <= (pair_idx+1)/2*4 + (pair_idx+1) mod 2;
                    bot_cpx  <= top_cpx + 2;
                    ram_addr <= cpx_to_addr(top_cpx, false);
                    st <= S1_RD_TOP_RE;
                end if;

            -- ==================== Stage-2 : distance 1 ====================
            when S2_RD_TOP_RE =>
                a_re <= wide_t(ram_din);
                ram_addr <= cpx_to_addr(top_cpx, true);
                st <= S2_RD_TOP_IM;

            when S2_RD_TOP_IM =>
                a_im <= wide_t(ram_din);
                ram_addr <= cpx_to_addr(bot_cpx, false);
                st <= S2_RD_BOT_RE;

            when S2_RD_BOT_RE =>
                b_re <= wide_t(ram_din);
                ram_addr <= cpx_to_addr(bot_cpx, true);
                st <= S2_RD_BOT_IM;

            when S2_RD_BOT_IM =>
                b_im <= wide_t(ram_din);
                k := tw_idx(2, pair_idx);             -- 0 1 2 3
                w_re <= TW_RE(k);
                w_im <= TW_IM(k);
                st <= S2_CALC;

            when S2_CALC =>
                -- 计算 a + b*Wk, a - b*Wk
                -- b' = b * Wk
                dn_re <= to_wide( mul_q15( signed(b_re(WIDTH-1 downto 0)), w_re) )
                       - to_wide( mul_q15( signed(b_im(WIDTH-1 downto 0)), w_im) );
                dn_im <= to_wide( mul_q15( signed(b_re(WIDTH-1 downto 0)), w_im) )
                       + to_wide( mul_q15( signed(b_im(WIDTH-1 downto 0)), w_re) );
                up_re <= a_re + dn_re;
                up_im <= a_im + dn_im;
                dn_re <= a_re - dn_re;
                dn_im <= a_im - dn_im;
                -- д�� Re
                ram_addr <= cpx_to_addr(top_cpx, false);
                ram_dout <= signed(up_re(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S2_WR_TOP_RE;

            when S2_WR_TOP_RE =>
                ram_addr <= cpx_to_addr(top_cpx, true);
                ram_dout <= signed(up_im(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S2_WR_TOP_IM;

            when S2_WR_TOP_IM =>
                ram_addr <= cpx_to_addr(bot_cpx, false);
                ram_dout <= signed(dn_re(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S2_WR_BOT_RE;

            when S2_WR_BOT_RE =>
                ram_addr <= cpx_to_addr(bot_cpx, true);
                ram_dout <= signed(dn_im(WIDTH-1 downto 0));
                ram_we   <= '1';
                st <= S2_WR_BOT_IM;

            when S2_WR_BOT_IM =>
                if pair_idx = 7 then          -- ȫ 8 �������
                    mag_idx  <= 0;
                    ram_addr <= cpx_to_addr(0, false);
                    st <= MAG_RD_RE;
                else
                    pair_idx <= pair_idx + 1;
                    top_cpx  <= pair_idx+1;
                    bot_cpx  <= top_cpx + 1;
                    ram_addr <= cpx_to_addr(top_cpx, false);
                    st <= S2_RD_TOP_RE;
                end if;

            -- ==================== ����ƽ�� ============================
            when MAG_RD_RE =>
                a_re <= wide_t(ram_din);                  -- Re
                ram_addr <= cpx_to_addr(mag_idx, true);   -- Im
                st <= MAG_RD_IM;

            when MAG_RD_IM =>
                a_im <= wide_t(ram_din);                  -- Im
                st <= MAG_CALC;

            when MAG_CALC =>
                mag32 := resize(a_re,34)*resize(a_re,34) +
                         resize(a_im,34)*resize(a_im,34);
                -- ���� 15 �� Q1.15
                ram_dout <= mag32(33 downto 18);
                ram_addr <= cpx_to_addr(mag_idx, false);  -- ����ԭ Re
                ram_we   <= '1';
                st <= MAG_WR;

            when MAG_WR =>
                if mag_idx = N-1 then
                    st <= DONE1;
                else
                    mag_idx <= mag_idx + 1;
                    ram_addr <= cpx_to_addr(mag_idx+1, false);
                    st <= MAG_RD_RE;
                end if;

            -- ==================== DONE ===============================
            when DONE1 =>
                done <= '1';
                if start='0' then
                    st <= IDLE;
                end if;

            end case;
        end if;
    end process;
end architecture;
